package TitanComms

    typedef enum [7:0] { 
        NOP = 0,
        WRITE = 1,
        READ = 2
     } instructions;

endpackage