package TitanComms;

    // typedef enum bit [7:0] { 
    //     NOP = 0,
    //     WRITE = 1,
    //     READ = 2
    //  } instructions;

    typedef enum int {
        NOP = 0, WRITE = 1, READ = 2
    } instructions;

endpackage